library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity squaretable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(7 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end squaretable;

architecture squaretable_arch of squaretable is
constant array_size 			: integer := 256 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal square_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;

begin  
  squaretable_proc: process(resetN, CLK)
    constant square_table : table_type := (
---start 0 v
X"3E80",
X"3D86",
X"3C8D",
X"3B97",
X"3AA3",
X"39B1",
X"38C1",
X"37D3",
X"36E7",
X"35FC",
X"3514",
X"342E",
X"3349",
X"3267",
X"3187",
X"30A8",
X"2FCC",
X"2EF1",
X"2E19",
X"2D42",
X"2C6E",
X"2B9B",
X"2ACA",
X"29FC",
X"292F",
X"2864",
X"279B",
X"26D5",
X"2610",
X"254D",
X"248C",
X"23CD",
X"2310",
X"2255",
X"219C",
X"20E5",
X"2030",
X"1F7D",
X"1ECB",
X"1E1C",
X"1D6F",
X"1CC4",
X"1C1B",
X"1B73",
X"1ACE",
X"1A2A",
X"1989",
X"18EA",
X"184C",
X"17B1",
X"1717",
X"1680",
X"15EA",
X"1556",
X"14C5",
X"1435",
X"13A7",
X"131B",
X"1292",
X"120A",
X"1184",
X"1100",
X"107E",
X"0FFE",
X"0F80",
X"0F04",
X"0E8A",
X"0E12",
X"0D9C",
X"0D28",
X"0CB6",
X"0C45",
X"0BD7",
X"0B6B",
X"0B01",
X"0A98",
X"0A32",
X"09CE",
X"096B",
X"090B",
X"08AC",
X"0850",
X"07F5",
X"079D",
X"0746",
X"06F1",
X"069F",
X"064E",
X"05FF",
X"05B2",
X"0568",
X"051F",
X"04D8",
X"0493",
X"0450",
X"040F",
X"03D0",
X"0393",
X"0358",
X"031F",
X"02E8",
X"02B3",
X"027F",
X"024E",
X"021F",
X"01F2",
X"01C6",
X"019D",
X"0176",
X"0150",
X"012D",
X"010B",
X"00EC",
X"00CE",
X"00B3",
X"0099",
X"0082",
X"006C",
X"0058",
X"0047",
X"0037",
X"0029",
X"001D",
X"0013",
X"000C",
X"0006",
X"0002",
X"0000",
X"0000",
X"0002",
X"0006",
X"000C",
X"0013",
X"001D",
X"0029",
X"0037",
X"0047",
X"0058",
X"006C",
X"0082",
X"0099",
X"00B3",
X"00CE",
X"00EC",
X"010B",
X"012D",
X"0150",
X"0176",
X"019D",
X"01C6",
X"01F2",
X"021F",
X"024E",
X"027F",
X"02B3",
X"02E8",
X"031F",
X"0358",
X"0393",
X"03D0",
X"040F",
X"0450",
X"0493",
X"04D8",
X"051F",
X"0568",
X"05B2",
X"05FF",
X"064E",
X"069F",
X"06F1",
X"0746",
X"079D",
X"07F5",
X"0850",
X"08AC",
X"090B",
X"096B",
X"09CE",
X"0A32",
X"0A98",
X"0B01",
X"0B6B",
X"0BD7",
X"0C45",
X"0CB6",
X"0D28",
X"0D9C",
X"0E12",
X"0E8A",
X"0F04",
X"0F80",
X"0FFE",
X"107E",
X"1100",
X"1184",
X"120A",
X"1292",
X"131B",
X"13A7",
X"1435",
X"14C5",
X"1556",
X"15EA",
X"1680",
X"1717",
X"17B1",
X"184C",
X"18EA",
X"1989",
X"1A2A",
X"1ACE",
X"1B73",
X"1C1B",
X"1CC4",
X"1D6F",
X"1E1C",
X"1ECB",
X"1F7D",
X"2030",
X"20E5",
X"219C",
X"2255",
X"2310",
X"23CD",
X"248C",
X"254D",
X"2610",
X"26D5",
X"279B",
X"2864",
X"292F",
X"29FC",
X"2ACA",
X"2B9B",
X"2C6E",
X"2D42",
X"2E19",
X"2EF1",
X"2FCC",
X"30A8",
X"3187",
X"3267",
X"3349",
X"342E",
X"3514",
X"35FC",
X"36E7",
X"37D3",
X"38C1",
X"39B1",
X"3AA3",
X"3B97",
X"3C8D",
X"3D86",
X"3E80"
 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= square_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end squaretable_arch;